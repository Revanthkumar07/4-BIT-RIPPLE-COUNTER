library verilog;
use verilog.vl_types.all;
entity RIPPER_vlg_vec_tst is
end RIPPER_vlg_vec_tst;
